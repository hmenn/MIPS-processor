module mips_testbench ();

endmodule
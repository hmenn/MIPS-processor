module mips_core(clock);
input clock;

endmodule

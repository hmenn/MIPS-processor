module mips_testbench ();
reg clock;
wire result;



endmodule
module mips_core();


endmodule
module alu_control_uni(ALUCtl,ALUOp,func);

  input [5:0]func;
  input [2:0]ALUOp;
  output [3:0] ALUCtl;




endmodule
